-- Instruction memory
-- May be implemented behaiorally using arrays

-- instructions are as follows:	
-- hex  -- instruction
-- 500A -- ldi $r0, 10
-- 5105 -- ldi $r1, 5
-- 5200 -- ldi $r2, 0
-- 5300 -- ldi $r3, 0
-- 5400 -- ldi $r4, 0
-- 5500 -- ldi $r5, 0
-- 5600 -- ldi $r6, 0
-- 5700 -- ldi $r7, 0
-- 0201 -- add $r2, $r0, $r1
-- 1301 -- mult $r3, $r0, $r1
-- 4401 -- sub $r4, $r0, $r1
-- 630B -- sh $r3, 0x0B
-- 640A -- sh $r4, 0x0A
-- 760A -- lh $r6, 0x0A
-- 770B -- lh $r7, 0x0B
